package sa_pkg;

endpackage
